module write_digit(
	input[3:0]a,
	input[3:0]b,
	input[3:0]c,
	input[3:0]d,
	input sa,
	input sb,
	input sc,
	input sd,
	output[6:0]a_to_g,
	output[3:0]en);
	
endmodule
